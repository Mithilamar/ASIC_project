interface tl_dll_intf(input logic clk);
endinterface
